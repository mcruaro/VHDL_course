--Implemente o trabalho 4 aqui. Envie pro Prof. somente esse arquivo no Logos