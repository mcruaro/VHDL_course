library IEEE;
use IEEE.std_Logic_1164.all;

package standards is

    --Constantes
    constant BUS_HIGH_INDEX  : integer := 7;

end standards;

