library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity senha is
    port (
        clock : in std_logic;
        reset : in std_logic;


    );
end senha;

architecture senha of senha is
    

    begin
       

end architecture;