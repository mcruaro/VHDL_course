--Implemente seu projeto aqui