library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity microondas is
    port (
        --Entrada
        clock : in std_logic;
        reset : in std_logic;
        --Entradas

        --Saidas
    );
end microondas;

architecture microondas of microondas is
    
    --Continuar
        
end architecture;